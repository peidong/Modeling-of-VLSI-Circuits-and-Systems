
VDD s 0 0
R1 s 1 2m
R2 1 2 2m
R3 2 3 3m
R4 2 n 3m
R5 n 5 4m
I1 1 0 3.408e-30
I2 2 0 6.592e-30
I3 3 0 1.6256e-29
I4 n 0 1.8418e-29
I5 5 0 1.0456e-29

.op
.print all
.plot all
.END
