* This is RC Circuit for hw 2
V1 6 0 DC=0V
R1 6 1 2m
R2 1 2 2m
R3 2 3 3m
R4 2 4 3m
R5 4 5 4m
I1 1 0 2n
I2 2 0 2n
I3 3 0 4n
I4 4 0 4n
I5 5 0 2n
.op
.end
