* This is RLC circuit
VDD 1 0 PULSE(0 1 0 10ps)
R1 4 5 2.916667e+00
R2 1 2 2.916667e+00
R3 7 8 2.916667e+00
C11 4 0 1.514721e-13
C12 6 0 1.514721e-13
C31 1 0 1.407739e-13
C32 3 0 1.407739e-13
C51 7 0 1.514721e-13
C52 9 0 1.514721e-13
C2 6 3 2.139635e-14
C4 9 3 2.139635e-14
L1 5 6 5.484192e-08
L2 2 3 5.484192e-08
L3 8 9 5.484192e-08
K1 L1 L2 7.389893e-01
K2 L1 L3 6.475001e-01
K3 L2 L3 7.389893e-01
.op
.TRAN 0.1ps 5ns
.print all
.plot all
.END
