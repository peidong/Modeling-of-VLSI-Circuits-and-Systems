* This is RC Circuit for hw 2
V1 6 0 DC=0V
R1 6 1 2m
R2 1 2 2m
R3 2 3 3m
R4 2 4 3m
R5 4 5 4m
I1 1 0 -2.20512e-40
I2 2 0 -4.27392e-40
I3 3 0 -10.49856e-40
I4 4 0 -12.01248e-40
I5 5 0 -6.84272e-40
.op
.end
