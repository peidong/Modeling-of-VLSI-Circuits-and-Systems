
VDD s 0 1
R1 s 1 2m
R2 1 2 2m
R3 2 3 3m
R4 2 n 3m
R5 n 5 4m
I1 1 0 0
I2 2 0 0
I3 3 0 0
I4 n 0 0
I5 5 0 0

.op
.print all
.plot all
.END
