*struct
V1 6 0 DC = 0V
R1 6 1 2m
R2 1 2 2m
R3 2 3 3m
R4 2 4 3m
R5 4 5 4m
I1 1 0 9.8e-29
I2 2 0 9.8e-29
I3 3 0 1.96e-28
I4 4 0 1.96e-28
I5 5 0 9.8e-29
.op
.end


